`timescale 1ns/1ps

`include "alu.v"
`include "calc.v" 
`include "decoder.v" 
`include "regfile.v"
`include "datapath.v"
`include "multicycle.v"
`include "ram.v"
`include "rom.v"
