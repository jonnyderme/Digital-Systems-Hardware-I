`timescale 1ns/1ps

//`include "calc_tb.v"
`include "multicycle_tb.v"
